package env_pkg;
   import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "decimal_encoding.sv"
  //`include "bfm.sv"
  `include "command_transaction.sv"
  `include "result_transaction.sv"
  `include "driver.sv"	
  `include "tester.sv"
  `include "command_monitor.sv"
  `include "coverage.sv"
  `include "result_monitor.sv"
  `include "scoreboard.sv"
  `include "env.sv"
  `include "random_test.sv"

endpackage 